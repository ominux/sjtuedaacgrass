inverter.cir -- a simple inverter
* The ideal opamp is modeled as a VCVS with a large gain.

R1 1 2 10k
R2 2 3 10k
E1 3 0 0 2 1e10
*E1 models the ideal opamp.

Vin 1 0 ac 1
.ac dec 10 1k 100k
.print ac V(3)
.end

