*bandgap.sp
.option post

****************************************
** Distributed RLC
****************************************

vin 1 0 dc 1 ac 1

r1 1 2 10k
c1 2 0 90.87n
r3 2 5 10k
r4 4 5 568.1k
c2 2 3 90.87n
r2 3 0 245.4
r5 4 0 10k
e1 5 0 3 4  1e+10

r6 5 6 10k
c3 6 0 44.37n
r7 6 9 9.558k
r8 8 9 17.45k
c4 6 7 44.37n
r9 7 0 9.774k
r10 8 0 10k
e2 9 0 7 8 1e+10 

r11 9 10 10k
c5 10 0 4.781n
r12 10 13 9.558k
r13 12 13 17.45k
c6 10 11 4.781n
r14 11 0 9.774k
r15 12 0 10k
e3 13 0 11 12 1e+10

.ac dec 100 100 10k
.print ac vm(13)

.end

