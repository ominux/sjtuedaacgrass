Self-Bias Inverter
VIN 20001 20002 ac 1
 
 

 
*netlist---------------------------------------
 

 
 
CL 20003 0 10p
 
M1 20003 20001 0 0 nch3 L=1u W=5u
rd_1 20003 20004 272.0000m
rs_1 0 20005 272.0000m
capbd_1 20004 0 4.7501f
capbs_1 20005 0 4.7501f
gm_1 20004 20005 20001 0 106.8048u
rds_1 20004 20005 5280857.10423
cgs_1 20001 20005 14.2486f
cgd_1 20001 20004 1.5789f
 
M2 20003 20001 0 0 pch3 L=1u W=10u
rd_2 20003 20006 144.0000m
rs_2 0 20007 144.0000m
capbd_2 20006 0 8.8966f
capbs_2 20007 0 8.8966f
gm_2 20006 20007 20001 0 73.5537u
rds_2 20006 20007 7126110.78252
cgs_2 20001 20007 34.1837f
cgd_2 20001 20006 2.7591f
 
M3 20008 20008 0 0 nch3 L=1u W=5u
rd_3 20008 20009 272.0000m
rs_3 0 20010 272.0000m
capbd_3 20009 0 4.7501f
capbs_3 20010 0 4.7501f
gm_3 20009 20010 20008 0 106.8048u
rds_3 20009 20010 5280857.10423
cgs_3 20008 20010 14.2486f
cgd_3 20008 20009 1.5789f
 
M4 20008 20008 0 0 pch3 L=1u W=10u
rd_4 20008 20011 144.0000m
rs_4 0 20012 144.0000m
capbd_4 20011 0 8.8966f
capbs_4 20012 0 8.8966f
gm_4 20011 20012 20008 0 73.5537u
rds_4 20011 20012 7126110.78252
cgs_4 20008 20012 34.1837f
cgd_4 20008 20011 2.7591f
 
E1 20002 0 20008 0 1
 
 
*extra control information---------------------
 

 
*.options post=2 nomod
 
.options list node post=2 probe
 
.op
 

 
*analysis--------------------------------------
 

 
.TRAN 1ns 300ns
 
*.DC VIN 0 5 0.1
 
.print ac VDB(20003) VP(20003)
 
*.ac dec 1000 1k 100g
 
.END
 

 
