Sallen-Key topology
vin 1 0 ac 1
r1 1 2 10k
r2 2 4 13k
c1 2 3 100p
c2 4 0 100p
e1 3 0 4 3 1e10
.print v(3)
.end
