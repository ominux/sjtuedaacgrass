Modified Sallen-Key topology
Vin 1 0 ac 1
R1 1 2 9.53k
R2 2 3 9.53k
C1 2 5 10n
C2 3 0 10n
Rf 5 4 3.65k
R0 4 0 10k
E1 5 0 3 4 1e10
.print v(5)
.end
