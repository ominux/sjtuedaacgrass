*bandgap.sp
.option post

****************************************
** Distributed RLC
****************************************

vin 1 0 dc 1
r1 1 2 50 
r2 3 4 50  
r3 5 6 50
r4 7 8 50
r5 9 10 50
r6 11 12 50
r7 13 14 50
r8 15 16 50
r9 17 18 50
r10 19 20 50
*r11 21 22 50
*r12 23 24 50
*r13 25 26 50
*r14 27 28 50
*r15 29 30 50
*r16 31 32 50
*r17 33 34 50
*r18 35 36 50
*r19 37 38 50
*r20 39 40 50
*r21 41 42 50
*r22 43 44 50
*r23 45 46 50
*r24 47 48 50
*r25 49 50 50
*r26 51 52 50
*r27 53 54 50
*r28 55 56 50
*r29 57 58 50
*r30 59 60 50
rload 19 0 100k 

c1 2 0 10p
c2 4 0 10p
c3 6 0 10p
c4 8 0 10p
c5 10 0 10p
c6 12 0 10p
c7 14 0 10p
c8 16 0 10p
c9 18 0 10p
c10 20 0 10p
*c11 22 0 10p
*c12 24 0 10p
*c13 26 0 10p
*c14 28 0 10p
*c15 30 0 10p
*c16 32 0 10p
*c17 34 0 10p
*c18 36 0 10p
*c19 38 0 10p
*c20 40 0 10p
*c21 42 0 10p
*c22 44 0 10p
*c23 46 0 10p
*c24 48 0 10p
*c25 50 0 10p
*c26 52 0 10p
*c27 54 0 10p
*c28 56 0 10p
*c29 58 0 10p
*c30 60 0 10p

l1 2 3 50n 
l2 4 5 50n  
l3 6 7 50n
l4 8 9 50n
l5 10 11 50n
l6 12 13 50n
l7 14 15 50n
l8 16 17 50n
l9 18 19 50n
l10 20 21 50n
*l11 22 23 50n
*l12 24 25 50n
*l13 26 27 50n
*l14 28 29 50n
*l15 30 31 50n
*l16 32 33 50n
*l17 34 35 50n
*l18 36 37 50n
*l19 38 39 50n
*l20 40 41 50n
*l21 42 43 50n
*l22 44 45 50n
*l23 46 47 50n
*l24 48 49 50n
*l25 50 51 50n
*l26 52 53 50n
*l27 54 55 50n
*l28 56 57 50n
*l29 58 59 50n
*l30 60 61 50n


.ac lin 1 100Meg
.print ac v(1,21)

.end

